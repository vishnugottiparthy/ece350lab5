// megafunction wizard: %LPM_DIVIDE%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_DIVIDE 

// ============================================================
// File Name: lpm_divider.v
// Megafunction Name(s):
// 			LPM_DIVIDE
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 17.0.2 Build 602 07/19/2017 SJ Lite Edition
// ************************************************************

//Copyright (C) 2017  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel MegaCore Function License Agreement, or other 
//applicable license agreement, including, without limitation, 
//that your use is for the sole purpose of programming logic 
//devices manufactured by Intel and sold by Intel or its 
//authorized distributors.  Please refer to the applicable 
//agreement for further details.

module lpm_divider (
	denom,
	numer,
	quotient,
	remain);

	input	[6:0]  denom;
	input	[7:0]  numer;
	output	[7:0]  quotient;
	output	[6:0]  remain;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: PRIVATE: PRIVATE_LPM_REMAINDERPOSITIVE STRING "TRUE"
// Retrieval info: PRIVATE: PRIVATE_MAXIMIZE_SPEED NUMERIC "-1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: USING_PIPELINE NUMERIC "0"
// Retrieval info: PRIVATE: VERSION_NUMBER NUMERIC "2"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_DREPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: LPM_HINT STRING "LPM_REMAINDERPOSITIVE=TRUE"
// Retrieval info: CONSTANT: LPM_NREPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_DIVIDE"
// Retrieval info: CONSTANT: LPM_WIDTHD NUMERIC "7"
// Retrieval info: CONSTANT: LPM_WIDTHN NUMERIC "8"
// Retrieval info: USED_PORT: denom 0 0 7 0 INPUT NODEFVAL "denom[6..0]"
// Retrieval info: USED_PORT: numer 0 0 8 0 INPUT NODEFVAL "numer[7..0]"
// Retrieval info: USED_PORT: quotient 0 0 8 0 OUTPUT NODEFVAL "quotient[7..0]"
// Retrieval info: USED_PORT: remain 0 0 7 0 OUTPUT NODEFVAL "remain[6..0]"
// Retrieval info: CONNECT: @denom 0 0 7 0 denom 0 0 7 0
// Retrieval info: CONNECT: @numer 0 0 8 0 numer 0 0 8 0
// Retrieval info: CONNECT: quotient 0 0 8 0 @quotient 0 0 8 0
// Retrieval info: CONNECT: remain 0 0 7 0 @remain 0 0 7 0
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_divider.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_divider.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_divider.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_divider.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_divider_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_divider_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
